library verilog;
use verilog.vl_types.all;
entity lab2_vlg_sample_tst is
    port(
        CLK             : in     vl_logic;
        input1          : in     vl_logic_vector(3 downto 0);
        input2          : in     vl_logic_vector(3 downto 0);
        reset           : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end lab2_vlg_sample_tst;
